module clocka(input clk,//ʱ������
				input sing_clk,
                 input clr,//�����ź�
                 input alarm_switch,//�л�Ϊ�趨����ģʽ
                 input set_button,//���ð�ť
                 input change_button,//�л���һ����ʾ��ť
                 input set_time_button,
                 output [0:6] r_s_g,//��ĸ�λ����ʾ
                 output [3:0] r_s,//���ʮλ����ʾ
                 output [3:0] r_m_g,//���ӵĸ�λ����ʾ
                 output [3:0] r_m,//���ӵ�ʮλ����ʾ
                 output [3:0] r_h_g,//Сʱ�ĸ�λ����ʾ
                 output [3:0] r_h,//Сʱ��ʮλ����ʾ
                 output reg speaker
                );//�����źź�����ź�
    parameter FREQ_C1 = 190;  // C1 Ƶ�� (262 Hz)
    parameter FREQ_D1 = 170;  // D1 Ƶ�� (294 Hz)
    parameter FREQ_E1 = 152;  // E1 Ƶ�� (330 Hz)
    parameter FREQ_F1 = 143;  // F1 Ƶ�� (349 Hz)
    parameter FREQ_G1 = 128;  // G1 Ƶ�� (392 Hz)
    parameter FREQ_A1 = 114;  // A1 Ƶ�� (440 Hz)
    parameter FREQ_B1 = 101;  // B1 Ƶ�� (494 Hz)
    parameter FREQ_C2 = 96;   // C2 Ƶ�� (523 Hz)
    reg [6:0] temp;
    reg [3:0] s_g, s, m_g, m, h_g, h; // ���ڴ洢��ǰʱ��ļĴ���
    reg [3:0] set_s_g, set_s, set_m_g, set_m, set_h_g, set_h; // �����������ӵļĴ���
    reg [2:0] set_pos; // ����λ�üĴ���
    reg sparkle;
    always@(posedge sing_clk)begin
	if((h_g==set_h_g&&h==set_h&&m_g==set_m_g&&m==set_m&&s==set_s&&set_time_button)||(m==4'b0000&&m_g==4'b0000))begin
	              if (temp == FREQ_C2-1) begin // ���������ӵ���ģ
                    speaker <= ~speaker; // ��ת����ź�
                    temp<= 0; // ����������
                end else 
                    temp = temp + 1; // �����������1
        end
        else
        speaker<=1'b0;
        end
    always @(posedge clk or negedge clr) begin//��ʱ���������ش���
        if(!clr) begin//�������־Ϊ1
            if(!alarm_switch) begin//�������־Ϊ0������ģʽΪ0
                h_g<=4'b0000;//Сʱ�ĸ�λ����
                h<=4'b0000;//Сʱ��ʮλ����
                m_g<=4'b0000;//���ӵĸ�λ����
                m<=4'b0000;//���ӵ�ʮλ����
                s_g<=4'b0000;//��ĸ�λ����
                s<=4'b0000;//���ʮλ����
            end
            else if(alarm_switch) begin//�������־Ϊ0������ģʽΪ1
                set_h_g<=4'b0000;//Сʱ�ĸ�λ����
                set_h<=4'b0000;//Сʱ��ʮλ����
                set_m_g<=4'b0000;//���ӵĸ�λ����
                set_m<=4'b0000;//���ӵ�ʮλ����
                set_s_g<=4'b0000;//��ĸ�λ����
                set_s<=4'b0000;//���ʮλ����
                set_pos<=3'b000;//����λ�üĴ�������
            end
        end
        else begin//�������־Ϊ1������ģʽΪ0
            if(s_g==4'b1001 && s==4'b0101) begin//����ǰ����Ϊ59
                s_g<=4'b0000;//��ĸ�λ����
                s<=4'b0000;//���ʮλ����
                if(m_g==4'b1001 && m==4'b0101) begin//����ǰ������Ϊ59
                    m_g<=4'b0000;//���ӵĸ�λ����
                    m<=4'b0000;//���ӵ�ʮλ����
                    if(h_g==4'b0011 && h==4'b0010) begin//����ǰСʱ��Ϊ23
                        h_g<=4'b0000;//Сʱ�ĸ�λ����
                        h<=4'b0000;//Сʱ��ʮλ����
                    end
                    else begin
                        if(h_g==4'b1001) begin//����ǰСʱ��Ϊ9
                            h_g<=4'b0000;//Сʱ�ĸ�λ����
                            h<=h+1;//Сʱ��ʮλ��һ
                        end
                        else begin//�������
                            h_g<=h_g+1;//Сʱ�ĸ�λ�ü�һ
                            h<=h;//Сʱ��ʮλ����
                        end
                    end
                end
                else begin//�������
                    if(m_g==4'b1001) begin//����ǰ������Ϊ9
                        m_g<=4'b0000;//���ӵĸ�λ����
                        m<=m+1;//���ӵ�ʮλ��һ
                    end
                    else begin//�������
                        m_g<=m_g+1;//���ӵĸ�λ�ü�һ
                        m<=m;//���ӵ�ʮλ����
                    end
                end
            end
            else if(s_g==4'b1001) begin//����λ����Ϊ9
                s_g<=4'b0000;//��λ����
                s<=s+1;//ʮλ��һ
            end
            else begin//��Ϊ�������
                s_g<=s_g+1;//��λ��һ
                s<=s;//ʮλ����
            end
            sparkle<=~sparkle;
            if(alarm_switch) begin
                if(change_button) begin//���л���һ����ʾ��ť
                    set_pos<=set_pos+1;//����λ�ü�һ
                    if(set_pos==3'b110)
                        set_pos<=3'b000;//������λ��Ϊ6������
                end
                if(set_button) begin//�����ð�ť����
                    case(set_pos)
                        3'b000: begin
                            if(set_s_g==4'b1001)//����ĸ�λΪ9������
                                set_s_g<=4'b0000;//��λ����
                            else
                            set_s_g<=set_s_g+1;//��ĸ�λ��һ
                        end
                        3'b001: begin
                            if(set_s==4'b0101)//�����ʮλΪ5������
                                set_s<=4'b0000;//ʮλ����
                            else
                            set_s<=set_s+1;//���ʮλ��һ
                        end
                        3'b010: begin
                            if(set_m_g==4'b1001)//�����ӵĸ�λΪ9������
                                set_m_g<=4'b0000;//��λ����
                            else
                              set_m_g<=set_m_g+1;//���ӵĸ�λ��һ
                        end
                        3'b011: begin
                            if(set_m==4'b0101)//�����ӵ�ʮλΪ5������
                                set_m<=4'b0000;//ʮλ����
                            else
                            set_m<=set_m+1;//���ӵ�ʮλ��һ
                        end
                        3'b100: begin
                            if(set_h_g==4'b0011)//��Сʱ�ĸ�λΪ3������
                                set_h_g<=4'b0000;//��λ����
                            else
                            set_h_g<=set_h_g+1;//���ӵ�ʮλ��һ
                        end
                        3'b101: begin
                            if(set_h==4'b0010)//��Сʱ��ʮλΪ2������
                                set_h<=4'b0000;//ʮλ����
                            else
                            set_h<=set_h+1;//Сʱ��ʮλ��һ
                        end
                    endcase
                end
                if(set_time_button)begin
				h_g<=set_h_g;//Сʱ�ĸ�λ����
                h<=set_h;//Сʱ��ʮλ����
                m_g<=set_m_g;//���ӵĸ�λ����
                m<=set_m;//���ӵ�ʮλ����
                s_g<=set_s_g;//��ĸ�λ����
                s<=set_s;//���ʮλ����
            end


            end
        end
        end
         assign   r_s_g= (alarm_switch) ? ((sparkle && set_pos==3'b000) ? turn_led(4'b1111) :turn_led(set_s_g) ) : turn_led(s_g);//��ĸ�λ����ʾ
         assign   r_s= (alarm_switch) ? ((sparkle && set_pos==3'b001) ? 4'b1111 : set_s) : s;//���ʮλ����ʾ
         assign   r_m_g= (alarm_switch) ? ((sparkle && set_pos==3'b010) ? 4'b1111 :set_m_g ): m_g;//���ӵĸ�λ����ʾ
         assign   r_m=(alarm_switch) ?((sparkle && set_pos==3'b011) ? 4'b1111 : set_m ) : m;//���ӵ�ʮλ����ʾ
         assign   r_h_g= (alarm_switch) ?((sparkle && set_pos==3'b100) ? 4'b1111 :set_h_g ): h_g;//Сʱ�ĸ�λ����ʾ
         assign   r_h=(alarm_switch) ?((sparkle && set_pos==3'b101) ? 4'b1111 : set_h) : h;//Сʱ��ʮλ����ʾ
    function[0:6] turn_led;
        input [3:0] g;
        begin
            case(g)
                4'b0000:
                    turn_led=7'b1111110;
                4'b0001:
                    turn_led=7'b0110000;
                4'b0010:
                    turn_led=7'b1101101;
                4'b0011:
                    turn_led=7'b1111001;
                4'b0100:
                    turn_led=7'b0110011;
                4'b0101:
                    turn_led=7'b1011011;
                4'b0110:
                    turn_led=7'b0011111;
                4'b0111:
                    turn_led=7'b1110000;
                4'b1000:
                    turn_led=7'b1111111;
                4'b1001:
                    turn_led=7'b1110011;
                default:
                    turn_led=7'b0000000;
            endcase
        end
    endfunction
endmodule
